module controller (
    input clk,
    input [53:0] decoded_instr
    
    
);

reg [4:0] states; //each bit stands for one state, one-hot coding
always @(posedge clk) 
begin
    
end




endmodule //controller