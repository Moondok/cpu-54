module instrument_decoder (
    input [31:0] raw_instruction,
    input ena,
    output reg[53:0] code
);
// here we translate mips 32 instrument to one hot code
wire [11:0] tmp={raw_instruction[31:26],raw_instruction[5:0]};

// we transform mips instruction into one-hot code to generate control signal
always @(*) 
begin
    if(ena)
    casex (tmp)
    //R-type
        12'b000000_100000: code<=54'b000000_00000000_00000000_00000000_00000000_00000000_00000001; //add
        12'b000000_100001: code<=54'b000000_00000000_00000000_00000000_00000000_00000000_00000010; //addu
        12'b000000_100010: code<=54'b000000_00000000_00000000_00000000_00000000_00000000_00000100; //sub
        12'b000000_100011: code<=54'b000000_00000000_00000000_00000000_00000000_00000000_00001000; //subu
        12'b000000_100100: code<=54'b000000_00000000_00000000_00000000_00000000_00000000_00010000; //and
        12'b000000_100101: code<=54'b000000_00000000_00000000_00000000_00000000_00000000_00100000; //or
        12'b000000_100110: code<=54'b000000_00000000_00000000_00000000_00000000_00000000_01000000; //xor
        12'b000000_100111: code<=54'b000000_00000000_00000000_00000000_00000000_00000000_10000000; //nor
        12'b000000_101010: code<=54'b000000_00000000_00000000_00000000_00000000_00000001_00000000; //slt
        12'b000000_101011: code<=54'b000000_00000000_00000000_00000000_00000000_00000010_00000000; //sltu
        12'b000000_000000: code<=54'b000000_00000000_00000000_00000000_00000000_00000100_00000000; //sll
        12'b000000_000010: code<=54'b000000_00000000_00000000_00000000_00000000_00001000_00000000; // srl
        12'b000000_000011: code<=54'b000000_00000000_00000000_00000000_00000000_00010000_00000000; // sra
        12'b000000_000100: code<=54'b000000_00000000_00000000_00000000_00000000_00100000_00000000; //sllv
        12'b000000_000110: code<=54'b000000_00000000_00000000_00000000_00000000_01000000_00000000; //srlv
        12'b000000_000111: code<=54'b000000_00000000_00000000_00000000_00000000_10000000_00000000; //srav
        12'b000000_001000: code<=54'b000000_00000000_00000000_00000000_00000001_00000000_00000000; //jr

        12'b001000_xxxxxx: code<=54'b000000_00000000_00000000_00000000_00000010_00000000_00000000; //addi
        12'b001001_xxxxxx: code<=54'b000000_00000000_00000000_00000000_00000100_00000000_00000000; //addiu
        12'b001100_xxxxxx: code<=54'b000000_00000000_00000000_00000000_00001000_00000000_00000000; //andi
        12'b001101_xxxxxx: code<=54'b000000_00000000_00000000_00000000_00010000_00000000_00000000; //ori
        12'b001110_xxxxxx: code<=54'b000000_00000000_00000000_00000000_00100000_00000000_00000000; //xori
        12'b001111_xxxxxx: code<=54'b000000_00000000_00000000_00000000_01000000_00000000_00000000; //lui
        12'b100011_xxxxxx: code<=54'b000000_00000000_00000000_00000000_10000000_00000000_00000000; //lw //23
        12'b101011_xxxxxx: code<=54'b000000_00000000_00000000_00000001_00000000_00000000_00000000; //sw //24
        12'b000100_xxxxxx: code<=54'b000000_00000000_00000000_00000010_00000000_00000000_00000000; //beq
        12'b000101_xxxxxx: code<=54'b000000_00000000_00000000_00000100_00000000_00000000_00000000;  //bne
        12'b001010_xxxxxx: code<=54'b000000_00000000_00000000_00001000_00000000_00000000_00000000; //slti
        12'b001011_xxxxxx: code<=54'b000000_00000000_00000000_00010000_00000000_00000000_00000000; //sltiu
        
        12'b000010_xxxxxx: code<=54'b000000_00000000_00000000_00100000_00000000_00000000_00000000; //j 
        12'b000011_xxxxxx: code<=54'b000000_00000000_00000000_01000000_00000000_00000000_00000000; //jal

        // new 23 instructions 
        12'b011100_100000: code<=54'b000000_00000000_00000000_10000000_00000000_00000000_00000000; // clz
        12'b000000_011011: code<=54'b000000_00000000_00000001_00000000_00000000_00000000_00000000; // divu
        12'b000000_011010: code<=54'b000000_00000000_00000010_00000000_00000000_00000000_00000000; // div 
        12'b011100_000010: code<=54'b000000_00000000_00000100_00000000_00000000_00000000_00000000; // mul 
        12'b000000_011001: code<=54'b000000_00000000_00001000_00000000_00000000_00000000_00000000; // mulu

        12'b000000_001001: code<=54'b000000_00000000_00010000_00000000_00000000_00000000_00000000; // jalr 
        12'b000001_xxxxxx: code<=54'b000000_00000000_00100000_00000000_00000000_00000000_00000000; // bgez
        12'b100001_xxxxxx: code<=54'b000000_00000000_01000000_00000000_00000000_00000000_00000000; // lh //38
        12'b100000_xxxxxx: code<=54'b000000_00000000_10000000_00000000_00000000_00000000_00000000; // lb //39
        12'b100100_xxxxxx: code<=54'b000000_00000001_00000000_00000000_00000000_00000000_00000000; // lbu//40 
        12'b100101_xxxxxx: code<=54'b000000_00000010_00000000_00000000_00000000_00000000_00000000; // lhu //41
        12'b101000_xxxxxx: code<=54'b000000_00000100_00000000_00000000_00000000_00000000_00000000; // sb 
        12'b101001_xxxxxx: code<=54'b000000_00001000_00000000_00000000_00000000_00000000_00000000; // sh

        12'b000000_010000: code<=54'b000000_01000000_00000000_00000000_00000000_00000000_00000000; // mfhi 
        12'b000000_010001: code<=54'b000000_10000000_00000000_00000000_00000000_00000000_00000000; // mthi 
        12'b000000_010010: code<=54'b000001_00000000_00000000_00000000_00000000_00000000_00000000; // mflo 
        12'b000000_010011: code<=54'b000010_00000000_00000000_00000000_00000000_00000000_00000000; // mtlo
        12'b010000_011000: code<=54'b000100_00000000_00000000_00000000_00000000_00000000_00000000; // eret
        12'b000000_001100: code<=54'b001000_00000000_00000000_00000000_00000000_00000000_00000000; // syscall 
        12'b000000_110100: code<=54'b010000_00000000_00000000_00000000_00000000_00000000_00000000; // teq
        12'b000000_001101: code<=54'b100000_00000000_00000000_00000000_00000000_00000000_00000000; //  break

        default: 
        begin
            if(raw_instruction[31:21]==11'b01000_000000)
                code<=54'b000000_00000000_00010000_00000000_00000000_00000000_00000000; // mfc0 44
            else if(raw_instruction[31:21]==11'b01000_000100)
                code<=54'b000000_00000000_00100000_00000000_00000000_00000000_00000000; // mtc0 45
            else
                code<=54'bz;
        end
            
    endcase
end
    


endmodule //instrument_decoder